/*

 #
 # This code is part of the research paper:
 # "Temporal Thermal Covert Channels in Cloud FPGAs"
 #
 # Copyright (C) Shanquan Tian, CASLAB @ Yale
 # Author: Shanquan Tian <shanquan.tian@yale.edu>
 #
 # MIT License
 #  
 # Permission is hereby granted, free of charge, to any person obtaining a copy of this software and associated 
 # documentation files (the ""Software""), to deal in the Software without restriction, including without limitation 
 # the rights to use, copy, modify, merge, publish, distribute, sublicense, and/or sell copies of the Software, and 
 # to permit persons to whom the Software is furnished to do so, subject to the following conditions:
 #  
 # The above copyright notice and this permission notice shall be included in all copies or substantial portions of the Software.
 #  
 # THE SOFTWARE IS PROVIDED *AS IS*, WITHOUT WARRANTY OF ANY KIND, EXPRESS OR IMPLIED, INCLUDING BUT NOT LIMITED TO THE 
 # WARRANTIES OF MERCHANTABILITY, FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE AUTHORS OR 
 # COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, 
 # ARISING FROM, OUT OF OR IN CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER DEALINGS IN THE SOFTWARE.
 # 

*/

module heater_1024(
    input enable,
    output wire [63:0] send
);

localparam HEATER_SIZE = 1024;

reg [10:0] heating_select = 0;
wire ro_heating_tick_selected;

mux_N_1  #( // HEATER_SIZE to 1 MUX
  .NWAY (HEATER_SIZE)
)
mux_heating (
  .select(heating_select),
  .ro_in(ro_heating_tick),
  .ro_selected(ro_heating_tick_selected)
);

reg ro_heating_reset = 0;

counter ro_heating_counter(
  .tick(ro_heating_tick_selected),
  .reset(ro_heating_reset),
  .val(send)
);


reg                   ro_heating_enable = 0;
wire[HEATER_SIZE-1:0] ro_heating_tick;

always @ (enable) begin
	ro_heating_enable = enable;
end

always @ (posedge enable) begin
    if (heating_select < HEATER_SIZE - 1) begin
    	heating_select <= heating_select + 1;
    end
	else begin
		heating_select <= 0;
	end
end



ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_0 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[0])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_1 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[1])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_2 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[2])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_3 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[3])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_4 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[4])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_5 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[5])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_6 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[6])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_7 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[7])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_8 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[8])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_9 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[9])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_10 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[10])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_11 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[11])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_12 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[12])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_13 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[13])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_14 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[14])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_15 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[15])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_16 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[16])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_17 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[17])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_18 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[18])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_19 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[19])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_20 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[20])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_21 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[21])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_22 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[22])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_23 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[23])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_24 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[24])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_25 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[25])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_26 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[26])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_27 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[27])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_28 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[28])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_29 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[29])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_30 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[30])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_31 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[31])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_32 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[32])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_33 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[33])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_34 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[34])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_35 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[35])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_36 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[36])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_37 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[37])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_38 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[38])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_39 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[39])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_40 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[40])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_41 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[41])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_42 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[42])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_43 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[43])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_44 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[44])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_45 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[45])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_46 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[46])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_47 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[47])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_48 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[48])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_49 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[49])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_50 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[50])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_51 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[51])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_52 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[52])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_53 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[53])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_54 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[54])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_55 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[55])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_56 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[56])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_57 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[57])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_58 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[58])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_59 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[59])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_60 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[60])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_61 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[61])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_62 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[62])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_63 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[63])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_64 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[64])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_65 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[65])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_66 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[66])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_67 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[67])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_68 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[68])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_69 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[69])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_70 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[70])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_71 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[71])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_72 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[72])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_73 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[73])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_74 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[74])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_75 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[75])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_76 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[76])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_77 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[77])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_78 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[78])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_79 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[79])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_80 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[80])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_81 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[81])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_82 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[82])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_83 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[83])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_84 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[84])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_85 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[85])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_86 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[86])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_87 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[87])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_88 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[88])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_89 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[89])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_90 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[90])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_91 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[91])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_92 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[92])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_93 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[93])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_94 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[94])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_95 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[95])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_96 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[96])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_97 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[97])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_98 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[98])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_99 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[99])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_100 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[100])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_101 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[101])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_102 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[102])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_103 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[103])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_104 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[104])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_105 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[105])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_106 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[106])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_107 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[107])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_108 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[108])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_109 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[109])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_110 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[110])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_111 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[111])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_112 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[112])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_113 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[113])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_114 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[114])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_115 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[115])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_116 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[116])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_117 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[117])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_118 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[118])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_119 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[119])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_120 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[120])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_121 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[121])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_122 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[122])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_123 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[123])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_124 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[124])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_125 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[125])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_126 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[126])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_127 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[127])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_128 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[128])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_129 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[129])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_130 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[130])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_131 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[131])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_132 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[132])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_133 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[133])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_134 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[134])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_135 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[135])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_136 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[136])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_137 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[137])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_138 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[138])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_139 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[139])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_140 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[140])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_141 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[141])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_142 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[142])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_143 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[143])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_144 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[144])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_145 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[145])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_146 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[146])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_147 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[147])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_148 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[148])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_149 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[149])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_150 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[150])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_151 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[151])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_152 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[152])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_153 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[153])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_154 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[154])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_155 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[155])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_156 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[156])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_157 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[157])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_158 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[158])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_159 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[159])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_160 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[160])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_161 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[161])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_162 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[162])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_163 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[163])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_164 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[164])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_165 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[165])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_166 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[166])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_167 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[167])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_168 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[168])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_169 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[169])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_170 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[170])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_171 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[171])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_172 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[172])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_173 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[173])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_174 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[174])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_175 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[175])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_176 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[176])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_177 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[177])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_178 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[178])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_179 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[179])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_180 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[180])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_181 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[181])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_182 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[182])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_183 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[183])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_184 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[184])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_185 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[185])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_186 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[186])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_187 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[187])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_188 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[188])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_189 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[189])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_190 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[190])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_191 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[191])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_192 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[192])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_193 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[193])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_194 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[194])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_195 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[195])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_196 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[196])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_197 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[197])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_198 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[198])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_199 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[199])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_200 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[200])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_201 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[201])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_202 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[202])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_203 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[203])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_204 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[204])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_205 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[205])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_206 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[206])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_207 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[207])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_208 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[208])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_209 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[209])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_210 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[210])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_211 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[211])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_212 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[212])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_213 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[213])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_214 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[214])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_215 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[215])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_216 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[216])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_217 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[217])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_218 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[218])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_219 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[219])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_220 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[220])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_221 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[221])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_222 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[222])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_223 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[223])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_224 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[224])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_225 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[225])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_226 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[226])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_227 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[227])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_228 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[228])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_229 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[229])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_230 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[230])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_231 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[231])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_232 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[232])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_233 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[233])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_234 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[234])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_235 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[235])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_236 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[236])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_237 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[237])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_238 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[238])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_239 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[239])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_240 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[240])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_241 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[241])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_242 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[242])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_243 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[243])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_244 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[244])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_245 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[245])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_246 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[246])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_247 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[247])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_248 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[248])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_249 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[249])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_250 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[250])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_251 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[251])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_252 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[252])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_253 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[253])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_254 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[254])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_255 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[255])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_256 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[256])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_257 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[257])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_258 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[258])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_259 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[259])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_260 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[260])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_261 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[261])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_262 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[262])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_263 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[263])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_264 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[264])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_265 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[265])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_266 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[266])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_267 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[267])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_268 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[268])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_269 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[269])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_270 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[270])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_271 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[271])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_272 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[272])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_273 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[273])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_274 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[274])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_275 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[275])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_276 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[276])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_277 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[277])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_278 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[278])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_279 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[279])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_280 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[280])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_281 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[281])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_282 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[282])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_283 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[283])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_284 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[284])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_285 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[285])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_286 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[286])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_287 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[287])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_288 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[288])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_289 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[289])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_290 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[290])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_291 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[291])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_292 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[292])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_293 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[293])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_294 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[294])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_295 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[295])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_296 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[296])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_297 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[297])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_298 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[298])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_299 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[299])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_300 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[300])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_301 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[301])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_302 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[302])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_303 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[303])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_304 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[304])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_305 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[305])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_306 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[306])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_307 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[307])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_308 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[308])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_309 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[309])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_310 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[310])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_311 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[311])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_312 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[312])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_313 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[313])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_314 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[314])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_315 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[315])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_316 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[316])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_317 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[317])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_318 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[318])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_319 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[319])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_320 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[320])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_321 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[321])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_322 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[322])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_323 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[323])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_324 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[324])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_325 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[325])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_326 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[326])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_327 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[327])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_328 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[328])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_329 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[329])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_330 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[330])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_331 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[331])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_332 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[332])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_333 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[333])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_334 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[334])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_335 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[335])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_336 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[336])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_337 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[337])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_338 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[338])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_339 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[339])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_340 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[340])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_341 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[341])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_342 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[342])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_343 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[343])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_344 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[344])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_345 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[345])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_346 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[346])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_347 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[347])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_348 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[348])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_349 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[349])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_350 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[350])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_351 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[351])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_352 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[352])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_353 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[353])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_354 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[354])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_355 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[355])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_356 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[356])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_357 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[357])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_358 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[358])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_359 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[359])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_360 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[360])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_361 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[361])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_362 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[362])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_363 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[363])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_364 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[364])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_365 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[365])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_366 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[366])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_367 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[367])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_368 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[368])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_369 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[369])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_370 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[370])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_371 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[371])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_372 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[372])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_373 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[373])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_374 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[374])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_375 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[375])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_376 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[376])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_377 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[377])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_378 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[378])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_379 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[379])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_380 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[380])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_381 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[381])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_382 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[382])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_383 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[383])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_384 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[384])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_385 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[385])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_386 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[386])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_387 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[387])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_388 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[388])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_389 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[389])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_390 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[390])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_391 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[391])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_392 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[392])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_393 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[393])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_394 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[394])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_395 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[395])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_396 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[396])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_397 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[397])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_398 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[398])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_399 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[399])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_400 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[400])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_401 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[401])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_402 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[402])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_403 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[403])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_404 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[404])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_405 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[405])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_406 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[406])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_407 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[407])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_408 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[408])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_409 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[409])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_410 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[410])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_411 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[411])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_412 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[412])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_413 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[413])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_414 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[414])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_415 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[415])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_416 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[416])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_417 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[417])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_418 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[418])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_419 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[419])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_420 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[420])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_421 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[421])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_422 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[422])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_423 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[423])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_424 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[424])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_425 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[425])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_426 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[426])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_427 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[427])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_428 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[428])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_429 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[429])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_430 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[430])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_431 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[431])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_432 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[432])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_433 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[433])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_434 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[434])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_435 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[435])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_436 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[436])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_437 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[437])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_438 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[438])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_439 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[439])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_440 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[440])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_441 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[441])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_442 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[442])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_443 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[443])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_444 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[444])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_445 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[445])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_446 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[446])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_447 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[447])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_448 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[448])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_449 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[449])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_450 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[450])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_451 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[451])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_452 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[452])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_453 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[453])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_454 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[454])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_455 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[455])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_456 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[456])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_457 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[457])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_458 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[458])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_459 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[459])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_460 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[460])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_461 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[461])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_462 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[462])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_463 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[463])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_464 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[464])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_465 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[465])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_466 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[466])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_467 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[467])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_468 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[468])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_469 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[469])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_470 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[470])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_471 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[471])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_472 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[472])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_473 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[473])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_474 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[474])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_475 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[475])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_476 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[476])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_477 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[477])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_478 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[478])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_479 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[479])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_480 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[480])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_481 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[481])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_482 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[482])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_483 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[483])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_484 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[484])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_485 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[485])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_486 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[486])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_487 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[487])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_488 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[488])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_489 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[489])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_490 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[490])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_491 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[491])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_492 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[492])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_493 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[493])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_494 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[494])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_495 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[495])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_496 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[496])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_497 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[497])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_498 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[498])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_499 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[499])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_500 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[500])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_501 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[501])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_502 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[502])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_503 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[503])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_504 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[504])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_505 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[505])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_506 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[506])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_507 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[507])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_508 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[508])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_509 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[509])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_510 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[510])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_511 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[511])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_512 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[512])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_513 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[513])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_514 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[514])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_515 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[515])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_516 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[516])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_517 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[517])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_518 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[518])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_519 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[519])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_520 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[520])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_521 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[521])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_522 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[522])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_523 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[523])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_524 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[524])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_525 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[525])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_526 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[526])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_527 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[527])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_528 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[528])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_529 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[529])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_530 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[530])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_531 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[531])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_532 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[532])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_533 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[533])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_534 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[534])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_535 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[535])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_536 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[536])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_537 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[537])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_538 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[538])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_539 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[539])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_540 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[540])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_541 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[541])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_542 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[542])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_543 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[543])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_544 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[544])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_545 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[545])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_546 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[546])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_547 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[547])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_548 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[548])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_549 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[549])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_550 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[550])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_551 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[551])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_552 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[552])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_553 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[553])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_554 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[554])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_555 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[555])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_556 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[556])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_557 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[557])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_558 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[558])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_559 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[559])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_560 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[560])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_561 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[561])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_562 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[562])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_563 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[563])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_564 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[564])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_565 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[565])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_566 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[566])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_567 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[567])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_568 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[568])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_569 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[569])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_570 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[570])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_571 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[571])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_572 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[572])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_573 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[573])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_574 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[574])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_575 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[575])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_576 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[576])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_577 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[577])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_578 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[578])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_579 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[579])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_580 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[580])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_581 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[581])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_582 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[582])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_583 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[583])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_584 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[584])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_585 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[585])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_586 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[586])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_587 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[587])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_588 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[588])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_589 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[589])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_590 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[590])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_591 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[591])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_592 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[592])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_593 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[593])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_594 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[594])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_595 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[595])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_596 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[596])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_597 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[597])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_598 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[598])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_599 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[599])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_600 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[600])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_601 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[601])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_602 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[602])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_603 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[603])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_604 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[604])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_605 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[605])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_606 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[606])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_607 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[607])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_608 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[608])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_609 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[609])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_610 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[610])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_611 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[611])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_612 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[612])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_613 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[613])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_614 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[614])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_615 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[615])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_616 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[616])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_617 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[617])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_618 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[618])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_619 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[619])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_620 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[620])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_621 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[621])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_622 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[622])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_623 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[623])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_624 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[624])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_625 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[625])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_626 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[626])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_627 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[627])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_628 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[628])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_629 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[629])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_630 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[630])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_631 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[631])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_632 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[632])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_633 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[633])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_634 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[634])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_635 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[635])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_636 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[636])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_637 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[637])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_638 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[638])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_639 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[639])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_640 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[640])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_641 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[641])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_642 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[642])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_643 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[643])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_644 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[644])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_645 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[645])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_646 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[646])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_647 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[647])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_648 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[648])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_649 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[649])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_650 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[650])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_651 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[651])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_652 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[652])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_653 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[653])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_654 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[654])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_655 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[655])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_656 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[656])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_657 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[657])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_658 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[658])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_659 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[659])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_660 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[660])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_661 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[661])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_662 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[662])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_663 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[663])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_664 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[664])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_665 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[665])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_666 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[666])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_667 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[667])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_668 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[668])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_669 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[669])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_670 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[670])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_671 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[671])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_672 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[672])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_673 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[673])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_674 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[674])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_675 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[675])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_676 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[676])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_677 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[677])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_678 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[678])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_679 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[679])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_680 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[680])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_681 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[681])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_682 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[682])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_683 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[683])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_684 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[684])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_685 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[685])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_686 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[686])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_687 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[687])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_688 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[688])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_689 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[689])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_690 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[690])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_691 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[691])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_692 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[692])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_693 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[693])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_694 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[694])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_695 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[695])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_696 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[696])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_697 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[697])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_698 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[698])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_699 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[699])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_700 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[700])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_701 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[701])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_702 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[702])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_703 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[703])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_704 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[704])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_705 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[705])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_706 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[706])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_707 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[707])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_708 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[708])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_709 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[709])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_710 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[710])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_711 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[711])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_712 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[712])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_713 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[713])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_714 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[714])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_715 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[715])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_716 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[716])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_717 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[717])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_718 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[718])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_719 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[719])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_720 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[720])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_721 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[721])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_722 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[722])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_723 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[723])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_724 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[724])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_725 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[725])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_726 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[726])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_727 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[727])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_728 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[728])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_729 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[729])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_730 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[730])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_731 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[731])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_732 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[732])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_733 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[733])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_734 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[734])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_735 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[735])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_736 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[736])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_737 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[737])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_738 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[738])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_739 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[739])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_740 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[740])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_741 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[741])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_742 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[742])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_743 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[743])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_744 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[744])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_745 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[745])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_746 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[746])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_747 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[747])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_748 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[748])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_749 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[749])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_750 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[750])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_751 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[751])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_752 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[752])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_753 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[753])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_754 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[754])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_755 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[755])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_756 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[756])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_757 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[757])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_758 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[758])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_759 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[759])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_760 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[760])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_761 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[761])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_762 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[762])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_763 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[763])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_764 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[764])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_765 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[765])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_766 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[766])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_767 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[767])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_768 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[768])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_769 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[769])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_770 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[770])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_771 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[771])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_772 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[772])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_773 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[773])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_774 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[774])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_775 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[775])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_776 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[776])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_777 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[777])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_778 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[778])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_779 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[779])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_780 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[780])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_781 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[781])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_782 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[782])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_783 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[783])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_784 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[784])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_785 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[785])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_786 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[786])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_787 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[787])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_788 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[788])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_789 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[789])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_790 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[790])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_791 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[791])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_792 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[792])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_793 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[793])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_794 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[794])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_795 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[795])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_796 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[796])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_797 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[797])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_798 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[798])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_799 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[799])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_800 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[800])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_801 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[801])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_802 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[802])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_803 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[803])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_804 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[804])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_805 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[805])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_806 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[806])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_807 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[807])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_808 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[808])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_809 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[809])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_810 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[810])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_811 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[811])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_812 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[812])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_813 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[813])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_814 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[814])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_815 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[815])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_816 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[816])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_817 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[817])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_818 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[818])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_819 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[819])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_820 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[820])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_821 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[821])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_822 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[822])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_823 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[823])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_824 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[824])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_825 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[825])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_826 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[826])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_827 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[827])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_828 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[828])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_829 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[829])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_830 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[830])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_831 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[831])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_832 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[832])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_833 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[833])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_834 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[834])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_835 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[835])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_836 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[836])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_837 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[837])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_838 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[838])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_839 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[839])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_840 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[840])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_841 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[841])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_842 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[842])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_843 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[843])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_844 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[844])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_845 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[845])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_846 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[846])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_847 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[847])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_848 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[848])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_849 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[849])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_850 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[850])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_851 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[851])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_852 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[852])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_853 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[853])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_854 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[854])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_855 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[855])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_856 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[856])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_857 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[857])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_858 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[858])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_859 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[859])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_860 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[860])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_861 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[861])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_862 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[862])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_863 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[863])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_864 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[864])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_865 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[865])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_866 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[866])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_867 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[867])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_868 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[868])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_869 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[869])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_870 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[870])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_871 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[871])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_872 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[872])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_873 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[873])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_874 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[874])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_875 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[875])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_876 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[876])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_877 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[877])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_878 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[878])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_879 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[879])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_880 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[880])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_881 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[881])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_882 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[882])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_883 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[883])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_884 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[884])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_885 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[885])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_886 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[886])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_887 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[887])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_888 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[888])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_889 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[889])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_890 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[890])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_891 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[891])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_892 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[892])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_893 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[893])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_894 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[894])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_895 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[895])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_896 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[896])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_897 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[897])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_898 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[898])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_899 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[899])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_900 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[900])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_901 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[901])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_902 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[902])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_903 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[903])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_904 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[904])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_905 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[905])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_906 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[906])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_907 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[907])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_908 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[908])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_909 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[909])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_910 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[910])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_911 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[911])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_912 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[912])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_913 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[913])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_914 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[914])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_915 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[915])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_916 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[916])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_917 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[917])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_918 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[918])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_919 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[919])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_920 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[920])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_921 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[921])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_922 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[922])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_923 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[923])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_924 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[924])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_925 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[925])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_926 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[926])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_927 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[927])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_928 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[928])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_929 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[929])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_930 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[930])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_931 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[931])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_932 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[932])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_933 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[933])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_934 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[934])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_935 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[935])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_936 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[936])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_937 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[937])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_938 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[938])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_939 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[939])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_940 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[940])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_941 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[941])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_942 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[942])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_943 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[943])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_944 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[944])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_945 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[945])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_946 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[946])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_947 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[947])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_948 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[948])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_949 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[949])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_950 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[950])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_951 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[951])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_952 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[952])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_953 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[953])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_954 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[954])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_955 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[955])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_956 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[956])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_957 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[957])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_958 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[958])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_959 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[959])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_960 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[960])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_961 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[961])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_962 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[962])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_963 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[963])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_964 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[964])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_965 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[965])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_966 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[966])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_967 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[967])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_968 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[968])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_969 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[969])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_970 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[970])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_971 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[971])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_972 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[972])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_973 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[973])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_974 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[974])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_975 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[975])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_976 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[976])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_977 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[977])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_978 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[978])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_979 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[979])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_980 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[980])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_981 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[981])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_982 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[982])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_983 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[983])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_984 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[984])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_985 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[985])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_986 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[986])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_987 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[987])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_988 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[988])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_989 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[989])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_990 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[990])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_991 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[991])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_992 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[992])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_993 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[993])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_994 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[994])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_995 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[995])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_996 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[996])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_997 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[997])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_998 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[998])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_999 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[999])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_1000 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[1000])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_1001 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[1001])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_1002 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[1002])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_1003 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[1003])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_1004 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[1004])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_1005 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[1005])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_1006 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[1006])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_1007 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[1007])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_1008 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[1008])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_1009 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[1009])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_1010 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[1010])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_1011 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[1011])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_1012 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[1012])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_1013 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[1013])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_1014 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[1014])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_1015 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[1015])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_1016 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[1016])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_1017 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[1017])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_1018 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[1018])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_1019 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[1019])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_1020 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[1020])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_1021 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[1021])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_1022 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[1022])
 );
ro_heater #(
  .RO_LENGTH (3)
)
ro_heating_1023 (
  .enable(ro_heating_enable),
  .out(ro_heating_tick[1023])
 );










endmodule
